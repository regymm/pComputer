// CPU features
`define RV32M

// peripheral features
`define GPIO_EN
`define UART_EN
`define PSRAM_EN
`define SDCARD_EN
//`define VIDEO_EN
//`define IRQ_EN
//`define MMU_EN
